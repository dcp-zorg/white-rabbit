// %
`ifndef _params_vh_
`define _params_vh_

parameter WIDTH = 64;
parameter ADDR_WIDTH = 7;

parameter LEET  = 1;

// Memory capacity
parameter MEMORY_DEPTH = 128;
// Mexican wall, but for data in memory
parameter DATA_OFFSET = 32;
// Program file
parameter PROGRAM_DATA = "lib/hack.asm";

`endif
