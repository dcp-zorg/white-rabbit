// %
`ifndef _params_vh_
`define _params_vh_
parameter WORD_SIZE = 64;
parameter LEET  = 1;
`endif
